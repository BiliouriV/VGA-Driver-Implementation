`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:36:51 11/27/2018 
// Design Name: 
// Module Name:    VRAM 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module VRAM(clk, reset, pixel_addr, haddr_enable, vaddr_enable, red_colour, green_colour, blue_colour);

input clk, reset;
input [13:0] pixel_addr;
input haddr_enable;
input vaddr_enable;

output red_colour;
output green_colour;
output blue_colour;

reg red_colour;
reg green_colour;
reg blue_colour;

wire red;
wire green;
wire blue;


//BLACK BACKGROUND VRAM --- FOR TESTING

  /* RAMB16_S1 #(
      .INIT(1'b0),  // Value of output RAM registers at startup
      .SRVAL(1'b0), // Output value upon SSR assertion
      .WRITE_MODE("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE

      // The forllowing INIT_xx declarations specify the initial contents of the RAM
      // Address 0 to 4095
      .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 4096 to 8191
      .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 8192 to 12287
      .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_23(256'h0000000000000000F0000000000000000000000000000000F000000000000000),
      .INIT_24(256'h0000000000000000F0000000000000000000000000000000F000000000000000),
      .INIT_25(256'h0000000000000000F0000000000000000000000000000000F000000000000000),
      .INIT_26(256'h0000000000000000F0000000000000000000000000000000F000000000000000),
      .INIT_27(256'h0000000000000000F0000000000000000000000000000000F000000000000000),
      .INIT_28(256'h0000000000000000F0000000000000000000000000000000F000000000000000),
      .INIT_29(256'h0000000000000000F0000000000000000000000000000000F000000000000000),
      .INIT_2A(256'h0000000000000000F0000000000000000000000000000000F000000000000000),
      .INIT_2B(256'h0000000000000000F0000000000000000000000000000000F000000000000000),
      .INIT_2C(256'h0000000000000000F0000000000000000000000000000000F000000000000000),
      .INIT_2D(256'h0000000000000000F0000000000000000000000000000000F000000000000000),
      .INIT_2E(256'h0000000000000000F0000000000000000000000000000000F000000000000000),
      .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 12288 to 16383
      .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
   ) RAMB16_S1_inst_blue (
      .DO(red_colour),      // 1-bit Data Output
      .ADDR(pixel_addr),  // 14-bit Address Input
      .CLK(clk),    // Clock
      .DI(1'b0),      // 1-bit Data Input
      .EN(1'b1),      // RAM Enable Input
      .SSR(1'b0),    // Synchronous Set/Reset Input
      .WE(1'b0)       // Write Enable Input
   );

  // End of RAMB16_S1_inst instantiation
						
						

/*green						
		
   // RAMB16_S1: 16kx1 Single-Port RAM
   //            Spartan-3
   // Xilinx HDL Language Template, version 14.6

   RAMB16_S1 #(
      .INIT(1'b0),  // Value of output RAM registers at startup
      .SRVAL(1'b0), // Output value upon SSR assertion
      .WRITE_MODE("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE

      // The forllowing INIT_xx declarations specify the initial contents of the RAM
      // Address 0 to 4095
      .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      // Address 4096 to 8191
      .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 8192 to 12287
      .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_23(256'h000000000000000F0000000000000000000000000000000F0000000000000000),
      .INIT_24(256'h000000000000000F0000000000000000000000000000000F0000000000000000),
      .INIT_25(256'h000000000000000F0000000000000000000000000000000F0000000000000000),
      .INIT_26(256'h000000000000000F0000000000000000000000000000000F0000000000000000),
      .INIT_27(256'h000000000000000F0000000000000000000000000000000F0000000000000000),
      .INIT_28(256'h000000000000000F0000000000000000000000000000000F0000000000000000),
      .INIT_29(256'h000000000000000F0000000000000000000000000000000F0000000000000000),
      .INIT_2A(256'h000000000000000F0000000000000000000000000000000F0000000000000000),
      .INIT_2B(256'h000000000000000F0000000000000000000000000000000F0000000000000000),
      .INIT_2C(256'h000000000000000F0000000000000000000000000000000F0000000000000000),
      .INIT_2D(256'h000000000000000F0000000000000000000000000000000F0000000000000000),
      .INIT_2E(256'h000000000000000F0000000000000000000000000000000F0000000000000000),
      .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 12288 to 16383
      .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
   ) RAMB16_S1_inst_green (
      .DO(green_colour),      // 1-bit Data Output
      .ADDR(pixel_addr),  // 14-bit Address Input
      .CLK(clk),    // Clock
      .DI(1'b0),      // 1-bit Data Input
      .EN(1'b1),      // RAM Enable Input
      .SSR(1'b0),    // Synchronous Set/Reset Input
      .WE(1'b0)       // Write Enable Input
   );

  // End of RAMB16_S1_inst instantiation
						
	
	
/*red

   // RAMB16_S1: 16kx1 Single-Port RAM
   //            Spartan-3
   // Xilinx HDL Language Template, version 14.6

   RAMB16_S1 #(
      .INIT(1'b0),  // Value of output RAM registers at startup
      .SRVAL(1'b0), // Output value upon SSR assertion
      .WRITE_MODE("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE

      // The forllowing INIT_xx declarations specify the initial contents of the RAM
      // Address 0 to 4095
      .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 4096 to 8191
      .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 8192 to 12287
      .INIT_20(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_23(256'h00000000000000F0000000000000000000000000000000F00000000000000000),
      .INIT_24(256'h00000000000000F0000000000000000000000000000000F00000000000000000),
      .INIT_25(256'h00000000000000F0000000000000000000000000000000F00000000000000000),
      .INIT_26(256'h00000000000000F0000000000000000000000000000000F00000000000000000),
      .INIT_27(256'h00000000000000F0000000000000000000000000000000F00000000000000000),
      .INIT_28(256'h00000000000000F0000000000000000000000000000000F00000000000000000),
      .INIT_29(256'h00000000000000F0000000000000000000000000000000F00000000000000000),
      .INIT_2A(256'h00000000000000F0000000000000000000000000000000F00000000000000000),
      .INIT_2B(256'h00000000000000F0000000000000000000000000000000F00000000000000000),
      .INIT_2C(256'h00000000000000F0000000000000000000000000000000F00000000000000000),
      .INIT_2D(256'h00000000000000F0000000000000000000000000000000F00000000000000000),
      .INIT_2E(256'h00000000000000F0000000000000000000000000000000F00000000000000000),
      .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 12288 to 16383
      .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
   ) RAMB16_S1_inst_red (
      .DO(blue_colour),      // 1-bit Data Output
      .ADDR(pixel_addr),  // 14-bit Address Input
      .CLK(clk),    // Clock
      .DI(1'b0),      // 1-bit Data Input
      .EN(1'b1),      // RAM Enable Input
      .SSR(1'b0),    // Synchronous Set/Reset Input
      .WE(1'b0)       // Write Enable Input
   );

*/

   // RAMB16_S1: 16kx1 Single-Port RAM
   //            Spartan-3
   // Xilinx HDL Language Template, version 14.7

		RAMB16_S1 #(
      .INIT(1'b0),  // Value of output RAM registers at startup
      .SRVAL(1'b0), // Output value upon SSR assertion
      .WRITE_MODE("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE

      // The forllowing INIT_xx declarations specify the initial contents of the RAM
      // Address 0 to 4095
      .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//red_white
      .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_red
      .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//red_white
      .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_red
      .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//red_white
      .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_red
      .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//red_white
      .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_red
      .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//green_white
      .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),		//white_green
      .INIT_0F(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//green_white
      // Address 4096 to 8191
      .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),		//white_green
      .INIT_12(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//green_white
      .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),		//white_green
      .INIT_15(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//green_white
      .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),		//white_green
      .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),		//white_blue
      .INIT_1A(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//blue_white
      .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),		//white_blue
      .INIT_1D(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//blue_white
      .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),		//white_blue
      // Address 8192 to 12287
      .INIT_20(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//blue_white
      .INIT_21(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_22(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),		//white_blue
      .INIT_23(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//blue_white
      .INIT_24(256'h000F0000F0000F0000F0000F0000F000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//black_white
      .INIT_25(256'h0FFF00FFF00FFF00FFF00FFF00FFF00F_0FFF00FFF00FFF00FFF00FFF00FFF00F),		//wwrgb_with white
      .INIT_26(256'h0FFF00FFF00FFF00FFF00FFF00FFF00F_000F0000F0000F0000F0000F0000F000),		//with white_with black
      .INIT_27(256'h000F0000F0000F0000F0000F0000F000_0FFF00FFF00FFF00FFF00FFF00FFF00F),		//with black_with white
      .INIT_28(256'h0FFF00FFF00FFF00FFF00FFF00FFF00F_0FFF00FFF00FFF00FFF00FFF00FFF00F),		//with white_with white
      .INIT_29(256'h0FFF00FFF00FFF00FFF00FFF00FFF00F_000F0000F0000F0000F0000F0000F000),		//with white_with black
      .INIT_2A(256'h000F0000F0000F0000F0000F0000F000_0FFF00FFF00FFF00FFF00FFF00FFF00F),		//with black_with white
      .INIT_2B(256'h0FFF00FFF00FFF00FFF00FFF00FFF00F_0FFF00FFF00FFF00FFF00FFF00FFF00F),		//with white_with white
      .INIT_2C(256'h0FFF00FFF00FFF00FFF00FFF00FFF00F_000F0000F0000F0000F0000F0000F000),		//with white_with black
      .INIT_2D(256'h000F0000F0000F0000F0000F0000F000_0FFF00FFF00FFF00FFF00FFF00FFF00F),		//with black_with white
      .INIT_2E(256'h0FFF00FFF00FFF00FFF00FFF00FFF00F_0FFF00FFF00FFF00FFF00FFF00FFF00F),		//with white_with white
      .INIT_2F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_000F0000F0000F0000F0000F0000F000),		//full white row_with black
      // Address 12288 to 16383
      .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),		
      .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),		
      .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),		
      .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),		
      .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),		
      .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
   ) RAMB16_RED_inst (
      .DO(red),      // 1-bit Data Output
      .ADDR(pixel_addr),  // 14-bit Address Input
      .CLK(clk),    // Clock
      .EN(1'b1),      // RAM Enable Input
      .SSR(reset),    // Synchronous Set/Reset Input
      .WE(1'b0)       // Write Enable Input
   );


		RAMB16_S1 #(
      .INIT(1'b0),  // Value of output RAM registers at startup
      .SRVAL(1'b0), // Output value upon SSR assertion
      .WRITE_MODE("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE

      // The forllowing INIT_xx declarations specify the initial contents of the RAM
      // Address 0 to 4095
      .INIT_00(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//red_white
      .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),		//white_red
      .INIT_03(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//red_white
      .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),		//white_red
      .INIT_06(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//red_white
      .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),		//white_red
      .INIT_09(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//red_white
      .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),		//white_red
      .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//green_white
      .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_green
      .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//green_white
      // Address 4096 to 8191
      .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_green
      .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//green_white
      .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_green
      .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//green_white
      .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_green
      .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),		//white_blue
      .INIT_1A(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//blue_white
      .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),		//white_blue
      .INIT_1D(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//blue_white
      .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),		//white_blue
      // Address 8192 to 12287
      .INIT_20(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//blue_white
      .INIT_21(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_22(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),		//white_blue
      .INIT_23(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//blue_white
      .INIT_24(256'h0000F0000F0000F0000F0000F0000F00_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//black_FULL white
      .INIT_25(256'h0FF0F0FF0F0FF0F0FF0F0FF0F0FF0F0F_0FF0F0FF0F0FF0F0FF0F0FF0F0FF0F0F),		//wwrgb_with white
      .INIT_26(256'h0FF0F0FF0F0FF0F0FF0F0FF0F0FF0F0F_0000F0000F0000F0000F0000F0000F00),		//with white_with black
      .INIT_27(256'h0000F0000F0000F0000F0000F0000F00_0FF0F0FF0F0FF0F0FF0F0FF0F0FF0F0F),		//with black_with white
      .INIT_28(256'h0FF0F0FF0F0FF0F0FF0F0FF0F0FF0F0F_0FF0F0FF0F0FF0F0FF0F0FF0F0FF0F0F),		//with white_with white
      .INIT_29(256'h0FF0F0FF0F0FF0F0FF0F0FF0F0FF0F0F_0000F0000F0000F0000F0000F0000F00),		//with white_with black
      .INIT_2A(256'h0000F0000F0000F0000F0000F0000F00_0FF0F0FF0F0FF0F0FF0F0FF0F0FF0F0F),		//with black_with white
      .INIT_2B(256'h0FF0F0FF0F0FF0F0FF0F0FF0F0FF0F0F_0FF0F0FF0F0FF0F0FF0F0FF0F0FF0F0F),		//with white_with white
      .INIT_2C(256'h0FF0F0FF0F0FF0F0FF0F0FF0F0FF0F0F_0000F0000F0000F0000F0000F0000F00),		//with white_with black
      .INIT_2D(256'h0000F0000F0000F0000F0000F0000F00_0FF0F0FF0F0FF0F0FF0F0FF0F0FF0F0F),		//with black_with white
      .INIT_2E(256'h0FF0F0FF0F0FF0F0FF0F0FF0F0FF0F0F_0FF0F0FF0F0FF0F0FF0F0FF0F0FF0F0F),		//with white_with white
      .INIT_2F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_0000F0000F0000F0000F0000F0000F00),		//full white row_with black
      // Address 12288 to 16383
      .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),		
      .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),		
      .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),		
      .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),		
      .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),		
      .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
   ) RAMB16_GREEN_inst (
      .DO(green),      // 1-bit Data Output
      .ADDR(pixel_addr),  // 14-bit Address Input
      .CLK(clk),    // Clock
      .EN(1'b1),      // RAM Enable Input
      .SSR(reset),    // Synchronous Set/Reset Input
      .WE(1'b0)       // Write Enable Input
   );


		RAMB16_S1 #(
      .INIT(1'b0),  // Value of output RAM registers at startup
      .SRVAL(1'b0), // Output value upon SSR assertion
      .WRITE_MODE("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE

      // The forllowing INIT_xx declarations specify the initial contents of the RAM
      // Address 0 to 4095
      .INIT_00(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//red_white
      .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),		//white_red
      .INIT_03(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//red_white
      .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),		//white_red
      .INIT_06(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//red_white
      .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),		//white_red
      .INIT_09(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//red_white
      .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),		//white_red
      .INIT_0C(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//green_white
      .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),		//white_green
      .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//green_white
      // Address 4096 to 8191
      .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),		//white_green
      .INIT_12(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//green_white
      .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),		//white_green
      .INIT_15(256'h00000000000000000000000000000000_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//green_white
      .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_00000000000000000000000000000000),		//white_green
      .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_blue
      .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//blue_white
      .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_blue
      .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//blue_white
      .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_blue
      // Address 8192 to 12287
      .INIT_20(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//blue_white
      .INIT_21(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_white
      .INIT_22(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//white_blue
      .INIT_23(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//blue_white
      .INIT_24(256'hF0000F0000F0000F0000F0000F0000F0_FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),		//black_FULL white
      .INIT_25(256'hFFF00FFF00FFF00FFF00FFF00FFF00FF_FFF00FFF00FFF00FFF00FFF00FFF00FF),		//wwrgb_with white
      .INIT_26(256'hFFF00FFF00FFF00FFF00FFF00FFF00FF_F0000F0000F0000F0000F0000F0000F0),		//with white_with black
      .INIT_27(256'hF0000F0000F0000F0000F0000F0000F0_FFF00FFF00FFF00FFF00FFF00FFF00FF),		//with black_with white
      .INIT_28(256'hFFF00FFF00FFF00FFF00FFF00FFF00FF_FFF00FFF00FFF00FFF00FFF00FFF00FF),		//with white_with white
      .INIT_29(256'hFFF00FFF00FFF00FFF00FFF00FFF00FF_F0000F0000F0000F0000F0000F0000F0),		//with white_with black
      .INIT_2A(256'hF0000F0000F0000F0000F0000F0000F0_FFF00FFF00FFF00FFF00FFF00FFF00FF),		//with black_with white
      .INIT_2B(256'hFFF00FFF00FFF00FFF00FFF00FFF00FF_FFF00FFF00FFF00FFF00FFF00FFF00FF),		//with white_with white
      .INIT_2C(256'hFFF00FFF00FFF00FFF00FFF00FFF00FF_F0000F0000F0000F0000F0000F0000F0),		//with white_with black
      .INIT_2D(256'hF0000F0000F0000F0000F0000F0000F0_FFF00FFF00FFF00FFF00FFF00FFF00FF),		//with black_with white
      .INIT_2E(256'hFFF00FFF00FFF00FFF00FFF00FFF00FF_FFF00FFF00FFF00FFF00FFF00FFF00FF),		//with white_with white
      .INIT_2F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF_F0000F0000F0000F0000F0000F0000F0),		//full white row_with black
      // Address 12288 to 16383
      .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),		
      .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),		
      .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),		
      .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),	
      .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),		
      .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),		
      .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
   ) RAMB16_BLUE_inst (
      .DO(blue),      // 1-bit Data Output
      .ADDR(pixel_addr),  // 14-bit Address Input
      .CLK(clk),    // Clock
      .EN(1'b1),      // RAM Enable Input
      .SSR(reset),    // Synchronous Set/Reset Input
      .WE(1'b0)       // Write Enable Input
   );


always @(posedge clk)
begin
	if (haddr_enable)
	begin
		if (vaddr_enable)
		begin
			red_colour = red;
			green_colour = green;
			blue_colour = blue;
		end
		else
		begin
			red_colour = 0;
			green_colour = 0;
			blue_colour = 0;
		end
	end
	else
	begin
		red_colour = 0;
		green_colour = 0;
		blue_colour = 0;
	end
end


endmodule
